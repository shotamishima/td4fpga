module data_selector(clk, rst, )
